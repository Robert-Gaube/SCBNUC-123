library verilog;
use verilog.vl_types.all;
entity count11_tb is
end count11_tb;
