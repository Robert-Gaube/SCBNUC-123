module seq3b (
  input [3:0] i,
  output reg o
);
  reg [3:0]var;
  reg [2:0]count;
  reg ultim;
  always@(*)
  begin
    var=i;
    ultim=i[0];
    count=3'b000;
    o=0;
    while(var>0)
    begin
      if(var[0]==ultim)
        count = count + 1;
      else
        count = 1;
      if(count==3)
        o=1;
      ultim=var[0];
      var=var/2;
    end
  end
endmodule

module seq3b_tb;
  reg [3:0] i;
  wire o;

  seq3b seq3b_i (.i(i), .o(o));

  integer k;
  initial begin
    $display("Time\ti\t\to");
    $monitor("%0t\t%b(%2d)\t%b", $time, i, i, o);
    i = 0;
    for (k = 1; k < 16; k = k + 1)
      #10 i = k;
  end
endmodule