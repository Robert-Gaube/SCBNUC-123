module main;
  initial
    $display("Ciao Lume!");
endmodule
    